library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity core is
	port (
		clk_in: in std_logic
	);
end core;


architecture rtl of core is
begin
end rtl;
