library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity bram is
	port(
		clka: in std_logic;
		ena: in std_logic;
		wea: in std_logic_vector(3 downto 0);
		addra: in std_logic_vector(11 downto 0);
		dia: in std_logic_vector(31 downto 0);
		doa: out std_logic_vector(31 downto 0);
		clkb: in std_logic;
		enb: in std_logic;
		addrb: in std_logic_vector(11 downto 0);
		dob: out std_logic_vector(31 downto 0)
	);
end bram;

architecture rtl of bram is
	type ram_type is array (0 to 4095) of std_logic_vector(31 downto 0);
	shared variable RAM: ram_type := (
X"008000ef", X"0000006f", X"000025b7", X"05800693", X"30858593", X"00b685b3", X"00000513", X"03200793",
X"06300713", X"00069603", X"00c787b3", X"0207d063", X"06478793", X"fe07cee3", X"0017b613", X"00268693",
X"00c50533", X"fed590e3", X"00008067", X"fef756e3", X"f9c78793", X"ff9ff06f", X"001c0011", X"ffe70008",
X"ffd00021", X"002a0002", X"fff60027", X"ffe6001d", X"002c0018", X"ffffffdb", X"0002fffc", X"fffaffd5",
X"001dffd4", X"ffd0002f", X"ffee000d", X"001e0012", X"0023ffd4", X"00020012", X"0032ffda", X"0012ffe4",
X"00200015", X"0012fff8", X"0018ffdf", X"fffa002e", X"0027fff7", X"00300007", X"ffe60029", X"0001ffcc",
X"ffd8ffff", X"0012ffc4", X"ffa9ffee", X"ffaa0049", X"0045ffd3", X"ffe1ffe8", X"fff4ffbb", X"0054ffb1",
X"00180053", X"ffb50046", X"ffdaffaf", X"001a0018", X"ffd0ffe6", X"fff6ffcc", X"0004ffa6", X"ffa80036",
X"fffd001f", X"ffbd005b", X"ffc30041", X"003fffe0", X"ffce0053", X"004bffa6", X"ffe9ffe6", X"ffc3ffe6",
X"ffbfffa7", X"003c00fa", X"ffd1028c", X"00320058", X"ff8fffc3", X"03370024", X"fcaf001a", X"001bffd2",
X"0029003a", X"ffd00044", X"000fffd6", X"0031ffea", X"0142004e", X"ffe4001c", X"ffdfffa1", X"ffe40038",
X"003f0025", X"fff8000d", X"0034ffc7", X"ffdcffc0", X"ffe4fff8", X"0031fec7", X"fff3ffa9", X"038f0018",
X"ff8bffdd", X"ffbf003c", X"fffd0022", X"00360034", X"fe8d0055", X"fff8ffbd", X"ffea029c", X"00330060",
X"ffc90008", X"001f0045", X"ffcf0053", X"00a5fd22", X"00550023", X"003cffd3", X"0020014c", X"ffe10024",
X"00e9ffea", X"0050fd42", X"0361ffe9", X"ffa2fffa", X"00120039", X"03bb00e1", X"ffd10022", X"ff9f0037",
X"0004fff7", X"002b003f", X"0012ffff", X"004b0007", X"ffb4ff20", X"004f000a", X"ffa5fc7e", X"fffdffd1",
X"0013ffb6", X"ffd30032", X"0036002e", X"001c0024", X"ffe50008", X"00290037", X"021cffd7", X"003a003c",
X"fffd004c", X"ffd3fcc1", X"ffb3ffb2", X"ffcefffe", X"fdc40018", X"ffa20003", X"ffcbfe03", X"022fffdd",
X"fedc0015", X"0010000a", X"032cff9e", X"000affd8", X"0010004a", X"005c00ff", X"ffb7029e", X"ffc50038",
X"fc56ffd7", X"ffacffc2", X"0059fffb", X"01a7ffe9", X"ff5e003e", X"fd46ffc7", X"002fffb0", X"fc7dfe63",
X"005cffbb", X"ff6f0142", X"0029003b", X"ffd90027", X"ffde0009", X"ffc6ffe4", X"ffc5022f", X"ffedffa7",
X"005efff3", X"004d0022", X"ffa5fffe", X"ffa2ffaa", X"ffc1ffbd", X"fffb01ae", X"00460005", X"ffbd001e",
X"ffe20043", X"ff7dffd9", X"0013ffeb", X"ffa00062", X"02620024", X"ffb80036", X"ffcfffa6", X"ffb3000b",
X"ffe2ffa3", X"004ffffb", X"003b0043", X"003fffe3", X"ffca0042", X"ff9bfdde", X"0004ffe4", X"0060fffa",
X"0143ffff", X"ffea01b3", X"ffb0ffb6", X"02920036", X"ffd20058", X"ffe90015", X"ffacffa7", X"00030048",
X"0028003c", X"ffcf0030", X"fffb0001", X"002eff3d", X"02aeffec", X"ffb00058", X"00510032", X"ffbdffe1",
X"fe72000f", X"fffffef3", X"fc2efd2e", X"ff670035", X"003d0027", X"02050007", X"ffedffe8", X"002d0013",
X"00460087", X"004303b6", X"fd60fef5", X"03800029", X"ffdfffbf", X"03730023", X"ffe5ffb8", X"ffafffaa",
X"ffa90051", X"0058000d", X"0034ffd0", X"ffccffd1", X"fd730075", X"ffa8ffdc", X"ffb9000c", X"00400019",
X"fff902ef", X"0256ffdf", X"0036ff9e", X"02fe001e", X"ffc4000f", X"ffff02b7", X"0027ffc8", X"ff9e0010",
X"00630065", X"fdccfeeb", X"ffeb0029", X"ffe9ffb1", X"00f60309", X"02330025", X"03100028", X"0038ffb0",
X"ffe1ffbb", X"00170003", X"ffa1feb5", X"003ffdcd", X"ffacfffb", X"0010ffd0", X"ffc10054", X"ffef004e",
X"ffe2ffc3", X"012d0003", X"0080001a", X"fff3fc24", X"0057fff2", X"0055000f", X"0030ffc3", X"0041fdb5",
X"003f0048", X"02ddfd0e", X"0248ffb1", X"0255ffaf", X"ffd8ffa2", X"ffa2ffbe", X"000f005e", X"0018fff1",
X"03270043", X"00560052", X"0014ffbe", X"005fffd7", X"0046001a", X"fffd01ae", X"ffd10003", X"fc86001f",
X"fff90201", X"0027003d", X"0376ffb5", X"0056ff9f", X"008c003c", X"0031ffa9", X"0017002e", X"000afffc",
X"ffc3feec", X"004c0018", X"ffd6ffc5", X"fff8fdee", X"fd480038", X"ffdaffad", X"0039fede", X"0063ffd9",
X"00370047", X"001cfe83", X"ffe6ffb5", X"004d0016", X"ffa2fffc", X"ffbc0044", X"000bff0a", X"ffcaffbf",
X"ffc6ffd2", X"ff9e0038", X"ffa2005e", X"001dfe53", X"00850363", X"00110029", X"fff7ffc6", X"fff40398",
X"ffe40001", X"0301ffb8", X"0012001f", X"00210052", X"fe890206", X"ff9effb2", X"fff0005c", X"001fffd4",
X"0041ffcd", X"ffef0028", X"fc910034", X"000e0003", X"001c017e", X"00170026", X"0365021b", X"ffe9ffd2",
X"fffdffa9", X"036e0316", X"ffd70233", X"0032ffbd", X"00370014", X"ffd1002a", X"ffb2ffd4", X"002cfd5d",
X"ffeafdbe", X"0015fccb", X"0012001c", X"002afd56", X"00080034", X"fc26ffbe", X"ffbdffb0", X"ffda0006",
X"ffdaffb0", X"ffe0ffab", X"005fffef", X"0019fffd", X"0013ffed", X"00b2ffc8", X"0037ffea", X"fc3afe9d",
X"fff8032a", X"ffc8fe7c", X"003301e5", X"ffceffe4", X"ffc0ffb1", X"ffccffe0", X"003dfebd", X"fdbdfebe",
X"01ddffdb", X"002e01fc", X"fda103cc", X"ffabfc69", X"0019fdf7", X"00200031", X"01dd0017", X"005c0047",
X"fe2cffca", X"fffb003b", X"feee0126", X"00410014", X"000d011f", X"ffb9fca8", X"0047fea8", X"ffc8004d",
X"014d005a", X"ffb10038", X"011e0004", X"ffb20059", X"003a0014", X"0336fec7", X"0005fffb", X"0052005c",
X"00290011", X"0032ffda", X"fc8effb9", X"004bffb5", X"ffd5012a", X"0005002d", X"004a0015", X"003affc9",
X"0279ffdc", X"002b0039", X"fff8000f", X"0178005d", X"0032fcf3", X"ffbc0037", X"ffef0038", X"0034ffb9",
X"004901b3", X"ffba0045", X"03520061", X"ffce002c", X"003efff8", X"fef00012", X"0055000f", X"00d6fff2",
X"ffd2002e", X"02efffcd", X"016b0025", X"ffaeffee", X"ffbc0120", X"fffdffa2", X"00520002", X"0020ffeb",
X"ffdb0052", X"ffdf0025", X"00340051", X"004a0033", X"ffcd004b", X"0034ffd4", X"0223002b", X"00b902f1",
X"0053004e", X"ffea0036", X"ffb90019", X"ffd1ffe0", X"002e003c", X"ffaf0050", X"037effdd", X"0045000e",
X"004affca", X"fffaffe8", X"fdcb0005", X"ffa3ffe2", X"001cfff9", X"ffd9ffab", X"003bffc1", X"fea7ffe2",
X"004bfd5e", X"fc74fe9e", X"000a026e", X"ffd00004", X"fffe0037", X"fffd0063", X"ffe1ffff", X"003cffca",
X"00540003", X"00e40028", X"ffa1005c", X"ffceff4f", X"003cffb9", X"001bffda", X"002f004b", X"000cff82",
X"0047011f", X"ffd9005f", X"01b9fff7", X"ff62ffa4", X"00050024", X"00330031", X"fe09036d", X"ffda00f1",
X"03cf004a", X"ffef0031", X"ffcb0013", X"001a0035", X"ffabffd7", X"01040016", X"ffedfff9", X"ffd0ffba",
X"0009010e", X"ffa80047", X"0057ffa9", X"000e0002", X"ffbd0054", X"ffdaffdf", X"ffdb004b", X"fff3000d",
X"ffff002b", X"00070033", X"ffe3003f", X"fdcd000f", X"ffed003a", X"feed0032", X"0047fff6", X"ffad002a",
X"ffc2ffec", X"ffe60058", X"ffffff9d", X"ffa1005d", X"ffc2ffdc", X"ffc3001d", X"0059002b", X"0041fff6",
X"0040030d", X"00100054", X"0013004c", X"fd260062", X"0399ffc1", X"fffc0053", X"ffacfff0", X"ffc7004d",
X"002e005b", X"fdde0059", X"00370011", X"ffe10033", X"ffc1ffa4", X"0010002f", X"00170014", X"0012ffd5",
X"ffdd0014", X"02960061", X"001a001c", X"ffeefff0", X"00040058", X"fffd001d", X"0084ffcb", X"ffdc0015",
X"005fffc5", X"ffba000f", X"0023ffb0", X"ffbe0042", X"001b003f", X"0044fe9a", X"01a7ffe9", X"ffe7003e",
X"ff2c003f", X"0032000c", X"0010ffe5", X"00240017", X"fff3ff9e", X"00340055", X"004efed2", X"ff3a018e",
X"ffce0060", X"0052ffd2", X"ffb0ff7f", X"0005fff3", X"ffa7ffb7", X"feb1ffc6", X"00580019", X"fff1ff5c",
X"005f003d", X"00010045", X"0110001e", X"ffb1ff23", X"001c00a5", X"0006002b", X"0052ffa0", X"fdba0052",
X"00520012", X"ffbafd83", X"fe29ffa3", X"ffd7fd87", X"ff040061", X"003f003b", X"0010ffda", X"003dffd7",
X"01510050", X"0045005e", X"0024ffc6", X"0053000f", X"003e039c", X"fff2ffd0", X"ffd5ffd8", X"0043002e",
X"ffecffdf", X"001c0017", X"0009fd1f", X"ffb3004d", X"00220035", X"ffbaffa9", X"00430046", X"03d3ffcf",
X"ffa2ffa9", X"fd43002d", X"003affee", X"ffd8003b", X"004c0051", X"004d00f3", X"fffb021c", X"000c0365",
X"00570385", X"fd800028", X"fdf60003", X"ffd1ff7a", X"ffca0036", X"ffed0374", X"000efef7", X"002b008f",
X"0013fd8b", X"004e0056", X"fff9ffd1", X"0037ffc5", X"fe6e000b", X"0109ffe3", X"ffc2ffa6", X"0063000b",
X"fcac0065", X"005cffd0", X"ffb70051", X"0001ffd7", X"ffc00037", X"ffe1ffec", X"ff40ff57", X"00600041",
X"005a0214", X"0021000f", X"001000ec", X"003f005e", X"00130002", X"003303b5", X"00060014", X"002dffb9",
X"fffe0348", X"029e005c", X"01aaffe6", X"ffc90012", X"fcde003f", X"005b0059", X"003cffbf", X"ffa10001",
X"fff8ff9f", X"ffed000f", X"004e003a", X"ffa7ffe0", X"ffd0001b", X"ffa50044", X"00cffd5f", X"fc19fffe",
X"fc1afffe", X"0042ffbe", X"001e0016", X"0053ffdd", X"ff6affa3", X"ffd90005", X"ffa8ffe9", X"0057ffe4",
X"0044fe29", X"ffadfe2c", X"ffabffef", X"0047ffd9", X"0053fc4d", X"0024ffdf", X"00190059", X"ffc70381",
X"0043ffd8", X"ffed02dd", X"0051fd0c", X"00350351", X"ffceffa7", X"ff1e0023", X"ffbc026a", X"fc4effae",
X"fffcfd1a", X"ff9effc6", X"0046000d", X"0055ffaf", X"fff6000f", X"002bffd7", X"00c203c8", X"0242002e",
X"ffc60016", X"0063fd05", X"fff60035", X"000effeb", X"001a0182", X"ffffffe7", X"ffa7fef2", X"004fffec",
X"ffab0042", X"ffff00ec", X"ffd30054", X"ffe90044", X"ffca0036", X"003ffff7", X"023effca", X"00be0006",
X"00baffba", X"ffbd0051", X"0079ff36", X"ffa2030d", X"fd29005e", X"ffb0fee8", X"00610057", X"ffbe0052",
X"01cd0057", X"ffdbfd07", X"002bfd78", X"003cff88", X"0053005f", X"0030ffd5", X"0019fffa", X"ffb7fff7",
X"ffb0fd1e", X"ffef0011", X"0002fff0", X"ffc3fff5", X"ffc503b1", X"0048fe6e", X"ffa60207", X"035bffdb",
X"005cffe6", X"ffc5000d", X"02c9fef2", X"0041ffac", X"ffca0023", X"00510036", X"ff14ff37", X"ffdf0059",
X"00520012", X"0141fff3", X"ff40fff8", X"004bfff8", X"00380019", X"fffb002c", X"01940370", X"00040011",
X"ffcdffcf", X"fff6000a", X"00320048", X"ff75fffd", X"03ceffb0", X"02ba003b", X"005a0029", X"ffcbfc85",
X"0055ffee", X"000dffb1", X"fddefd95", X"03260047", X"ffec0045", X"ffaaffb0", X"00510005", X"0040ffc0",
X"0058000c", X"0011feb5", X"0021fffd", X"00150117", X"fff9fd6d", X"004bffe7", X"004b02dc", X"000901ed",
X"0072fd81", X"0052ffac", X"ff790206", X"005affae", X"fd2c01e2", X"ffe10007", X"fff4ffd2", X"0021005c",
X"00bdffd8", X"fd16004d", X"019c0022", X"03bafff7", X"fffdfc4f", X"002bffd8", X"00500014", X"0006ffaf",
X"fe500010", X"fffafff7", X"ffa8ffa2", X"ffbbffd5", X"03a2005b", X"fd8f001d", X"0049ff9e", X"0014ffaa",
X"0009022d", X"0028ffc9", X"ffd6000f", X"003f002a", X"00390044", X"001a003a", X"ffc4ffa3", X"00060005",
X"ffbcffdd", X"ffa9ffe5", X"ffaf0036", X"ff7e000e", X"028afff1", X"ffea005f", X"ffb1feea", X"0040febf",
X"00600024", X"0005ffd2", X"003effc5", X"0052002a", X"0131000d", X"ffdaffc2", X"0055000f", X"ff54000f",
X"fffcff7f", X"ffc2005a", X"ffadffda", X"ffabffe0", X"ffa70059", X"fff303c3", X"00410055", X"ffd5ff9e",
X"fd090048", X"00030034", X"003bfc31", X"ffb1fff5", X"005aff23", X"0051001d", X"0292ffed", X"001c0047",
X"ffd3ffda", X"ff3b002d", X"fff60007", X"03790060", X"02cdffab", X"ffb4003b", X"0003031d", X"0018ffe8",
X"0131ffe8", X"ffd20041", X"ffb3fd91", X"ffe301ad", X"ff7d000d", X"000effae", X"010affab", X"ffaeffcb",
X"fff90038", X"0215005b", X"ffd30043", X"ffa4ffb5", X"fffb0067", X"0013000e", X"fe67005a", X"ffda03aa",
X"0048003a", X"00490039", X"ffc90030", X"00220015", X"035cffcc", X"fc74fff8", X"ffacffc0", X"000bffcc",
X"fff7004d", X"ff9f0015", X"ffda0061", X"fc2b0026", X"0055ffc8", X"ffd6fffa", X"001dff19", X"0059ffa8",
X"01780001", X"001b0018", X"0056ffe5", X"0040000e", X"00010060", X"001f0027", X"0041fff7", X"ffa1ffa5",
X"0284fc7b", X"00090038", X"ffef0008", X"00090015", X"005b004f", X"003efedf", X"00150047", X"fd310023",
X"02550016", X"0056fff5", X"00490058", X"00200020", X"0052ffac", X"00030002", X"fff40009", X"0016ffe0",
X"ffcbffa6", X"ffef0035", X"002affad", X"ffb8001e", X"fc580026", X"026dfe0a", X"0041ffe7", X"038803a7",
X"ffa6005a", X"ffd1ffcb", X"0027ffed", X"022dffd7", X"001affc2", X"ffe9013c", X"0027ffe0", X"fff100d7",
X"0017ffd3", X"ffd10021", X"fff0ffb2", X"fc500014", X"ffed0036", X"ffe70013", X"ffccffe9", X"0035015b",
X"025b0060", X"ffecff9d", X"005703e7", X"fffeffbe", X"004c0017", X"fffc0003", X"fdcb0045", X"02e90029",
X"0042fcac", X"01f7fffe", X"fc220063", X"0136005a", X"005efffb", X"0006ffdc", X"003dfda3", X"025fffe6",
X"0002ffa3", X"fc6d03d9", X"fd45000f", X"0053ffff", X"fed8ffa9", X"00330031", X"fe950045", X"001cfd22",
X"ffdd0008", X"000cfdd4", X"027bffe3", X"0001ffdc", X"ff9e002e", X"ffe50034", X"0046fd7d", X"001802e3",
X"fc41fffc", X"001e01d6", X"ffcaffd2", X"004fffd4", X"0043fde9", X"ffd502a4", X"ffa60062", X"002cfff8",
X"ffa4ffcc", X"ffa5fce1", X"fffefd9e", X"00340002", X"007b002d", X"0042ffec", X"00430043", X"03b2005a",
X"0027005b", X"00410045", X"003dffcd", X"ffc8002e", X"ffa80058", X"fffbffe1", X"00d4ffb4", X"ffc3fe49",
X"00010063", X"ffd9ffcf", X"ffcbffca", X"fd680046", X"003d0239", X"0044fff7", X"00130051", X"ffc20062",
X"0033ffce", X"ffd5fff6", X"ffcd01e5", X"ff0a0052", X"ffabfdd6", X"0035000e", X"ffff002f", X"ffbe0048",
X"005f0042", X"ffae0057", X"fff7ffbc", X"fe890046", X"002d0025", X"02890033", X"ffe9005a", X"fd84ffe1",
X"00140050", X"ff31ffa3", X"0020ffe0", X"ffeaffaf", X"ffa80003", X"004fffea", X"ff94001f", X"01540008",
X"008dffaf", X"001b0049", X"005b0135", X"ff90ffa8", X"0053004f", X"fe2b0133", X"005502cb", X"ffe7003f",
X"ffb40009", X"0038fceb", X"fef2ffda", X"ffe9fff9", X"ffc4ff9f", X"001fffd5", X"0048ffe1", X"ffd903c7",
X"ffe90062", X"ffb60039", X"00610062", X"000c02eb", X"ffbc0038", X"ffc3003d", X"0212ffcf", X"ffcf0042",
X"0024ff9e", X"001f0040", X"03530012", X"004dffb3", X"ffe800d4", X"000bffa8", X"fcb90008", X"ffb2ffee",
X"0016ffac", X"0038ffea", X"002fffc8", X"0048ffd1", X"ffacffb8", X"ffd2ffba", X"00120015", X"ffc4feeb",
X"ffe9fffe", X"ffe4001d", X"ffedffb2", X"ffba0016", X"03e40047", X"000e0056", X"004a001a", X"004f0015",
X"fff3ffc7", X"ffd4ffce", X"000f0040", X"ffe0ff8d", X"ff75ffe5", X"ffc2fc7a", X"0038ffaf", X"004d0004",
X"ffaf003c", X"005effb7", X"ffdbffa2", X"004500e5", X"ffcbffe7", X"023effad", X"ffe10359", X"fdc3ff81",
X"005c01fc", X"fd72fd16", X"000cffcd", X"ffdc004b", X"01360300", X"0055001e", X"fcb1ffd2", X"ffc2ffb0",
X"0137002a", X"03190103", X"0051ffd2", X"02eb0021", X"ffb501a6", X"0006004b", X"0029fffa", X"ffa4fc4b",
X"0044ff9b", X"001cffb5", X"ffca01d1", X"ff9f0042", X"0032ffc9", X"ffa8026f", X"ffa2fc58", X"fdc6ffdd",
X"ffc30005", X"003e0043", X"0038ffdc", X"002bffa8", X"ffaf000b", X"ffecffd1", X"0010fe06", X"02d7fff0",
X"ffdeffc9", X"ffb8fcb8", X"fff9ffed", X"ffa00060", X"0017ffe9", X"ffa20036", X"ffe4ffa2", X"fffbffd0",
X"000bfff8", X"ffecffa8", X"0012026c", X"0010ffde", X"00600068", X"00360026", X"fff90198", X"ffecffe8",
X"ffb8005b", X"ffcd0373", X"ff52003f", X"0008ffa7", X"01befff8", X"ffaf0044", X"fe6fffd2", X"fff7ffb3",
X"ffe6ffaa", X"004dfce8", X"033500a3", X"005bfcb0", X"003cfd7e", X"ffad001d", X"fe060047", X"ffb4ffcb",
X"ff72005d", X"fffafc49", X"000fffa5", X"ffa1004d", X"fcf80048", X"ffc2ffa0", X"0352ffc9", X"ffc0ffb8",
X"fffe0003", X"005d0002", X"ffbc0027", X"00080024", X"ffdfffc7", X"fe230052", X"01b5004d", X"ffa2003f",
X"0002003b", X"ffdeffd8", X"ffe7ffbf", X"00490061", X"ffff001b", X"ffacfff2", X"004b02d4", X"005bffa5",
X"ffc1016b", X"ffe30129", X"01ffffb1", X"0022016e", X"001b0022", X"0031003c", X"0112fe8e", X"ff840032",
X"0005fffb", X"0005fffb", X"ffd2005b", X"ffa8ffc7", X"ffe2feae", X"0042fffa", X"001f004d", X"ffc7ffd5",
X"004f0012", X"ffde0005", X"0226ffbc", X"003300c7", X"ffa101ef", X"ffcd004a", X"001fffe9", X"ff9dffad",
X"ffcf02d3", X"ffe4ffb9", X"004cff84", X"0060ffb8", X"0244ffee", X"ffdfff9d", X"00410046", X"004affd9",
X"fe2affa5", X"00410060", X"ffb0ffec", X"ffafffed", X"001dffdc", X"005affa3", X"001d002c", X"001c00d1",
X"ffff0003", X"ff95ffd3", X"0060ffdf", X"0008000e", X"ffd50109", X"ffe8ffdf", X"00020062", X"fe650219",
X"ffa3004d", X"feb40122", X"000c0014", X"0374ffac", X"fd3effd9", X"00100008", X"0017ffb1", X"fd28ffe9",
X"0005ffb8", X"ff9ffffb", X"ffde0033", X"0039ffec", X"0131ffc2", X"0005ffcd", X"fff2fe10", X"028e0028",
X"0047ffda", X"0012ffa7", X"001100b7", X"0004ffbe", X"ffb5003e", X"003c000f", X"004f0015", X"ffb70020",
X"0034fff9", X"fff8fec7", X"fcabfffa", X"ffeffff9", X"ffb80048", X"ffcefff2", X"ffa50033", X"0012005b",
X"ffa3fff4", X"ffdcffc0", X"0024ffe9", X"ffe6fff3", X"fffbffc2", X"fc510125", X"0011ffce", X"005f004f",
X"0056ffeb", X"0008ff05", X"016affae", X"003c0003", X"0030ffc1", X"000b0001", X"ffccffc4", X"ffadff1b",
X"ffb1002b", X"fffbffec", X"039fffb5", X"ffaeffe5", X"fff2010a", X"003f001e", X"00abffde", X"ffbcffe0",
X"0007005d", X"00b1fff4", X"0015ffaa", X"ffbbffe1", X"ffabfec2", X"0046ffb9", X"ffde0048", X"0050ff9f",
X"0009ff8b", X"0063005b", X"ffc0ff9d", X"ffcd004a", X"004fffc4", X"0332ffd6", X"0266ffca", X"ffedfd49",
X"ffddfc2d", X"ffcdfe1a", X"ffe40051", X"0013ffa4", X"000dffe3", X"000cffae", X"ffa10063", X"01250035",
X"0026ffa1", X"fed2ffcb", X"000a0013", X"002fffc7", X"004a0019", X"ffbf0035", X"ffd7000d", X"ffbdffbc",
X"ffe7ffba", X"ffa6ffce", X"02fbffa7", X"ffd0035f", X"0052ffbd", X"ff9effc6", X"ffa1fde7", X"002d0025",
X"ffe602cc", X"fee9ff9e", X"ffc5ffbe", X"ffe8ffb5", X"001e01a8", X"ffd3000f", X"ffb3ffba", X"0019fe9f",
X"ffc80023", X"ffcf0060", X"0015fd11", X"ffd5002f", X"ffc6ffbd", X"001f0048", X"0036ffaa", X"0364001d",
X"0019ffbc", X"002a005a", X"00590036", X"ffb7ffe5", X"019c0021", X"ffa9003e", X"0016ffd1", X"ffbeffcb",
X"ffb70060", X"ff9d0001", X"03100014", X"000d031b", X"fd3cfd9b", X"0045ffc3", X"00530011", X"fddeffca",
X"0321031f", X"ffe1ffac", X"ffeaffb2", X"ffd50059", X"003b004a", X"fc71ffc0", X"000b0035", X"000b015b",
X"0044000e", X"ffe10007", X"fe0bffbb", X"0063ff9e", X"fe7cffab", X"00080028", X"00050185", X"03670041",
X"ffc3fce2", X"001a0036", X"002fffe6", X"005fffdf", X"0324ffad", X"03b4001a", X"0005fff7", X"fff4004b",
X"ffd3ffee", X"0009ffee", X"010a0009", X"00370022", X"ffa20053", X"ff470029", X"ffb6ffd1", X"005bffb1",
X"ffacfff9", X"fc3cffdc", X"fdde002e", X"0009fff7", X"00280059", X"ffcbffff", X"0046fe25", X"ffc2fff8",
X"003c0028", X"005b003c", X"ffcb0031", X"00130022", X"0038fff6", X"ffdeffce", X"ffa4021a", X"000cfc74",
X"ffa6fff4", X"00030058", X"00380002", X"0006ffbf", X"013dffbf", X"fff9ff68", X"ffc40007", X"00190038",
X"002ffc20", X"0030fff3", X"fd70ffcc", X"fd0f000f", X"02bd0039", X"ffd30052", X"001301d3", X"ffe80036",
X"ffdb0020", X"001ffffe", X"005b003d", X"003afdf7", X"0059ff0e", X"ffd2005a", X"004d0398", X"0005ffb3",
X"ffa90052", X"fff0fe6c", X"ffd0ffd4", X"01a00070", X"fff9ff28", X"020afffa", X"ffe7005b", X"ffdafe4b",
X"ffb6fc84", X"ffe1fd86", X"ffc10024", X"00280012", X"01f8fffc", X"ffd80028", X"03090003", X"004bfe39",
X"fffc0057", X"003affad", X"ffbbfd15", X"0013003a", X"fff60051", X"ffbeffa6", X"fffeffce", X"0007ffae",
X"fe92fff9", X"ffdb0362", X"ffa6001b", X"ff360002", X"038a004f", X"001ffff0", X"0040ffcc", X"0024ffac",
X"ffd802c6", X"0016ffed", X"0039fd9d", X"0040ffcb", X"fff8000e", X"004c0006", X"0021024d", X"02ec0030",
X"0060fff5", X"000cffab", X"ffa2ffd2", X"00370046", X"00430111", X"00570371", X"fffffffc", X"ffa6ff9f",
X"00040057", X"ffc20060", X"ffb2003e", X"0001001c", X"00d8ffbd", X"0013ffed", X"004b0027", X"0061fd36",
X"ff9d0003", X"fff8ffa0", X"002ffe0d", X"0029ffc7", X"0021ffb7", X"0001000e", X"003fffd3", X"ffd1ffaa",
X"005b0014", X"00660062", X"ffea0057", X"00560024", X"ff2d0018", X"002cff27", X"002a001e", X"00c7ff9e",
X"0022ffde", X"005a0032", X"ffe0001c", X"ffc70040", X"0069001b", X"ffea002f", X"012dffdd", X"ffefffcf",
X"fcf6ffea", X"0006fda2", X"02c4ffe7", X"ffb10024", X"ffe10004", X"ffa4fff3", X"00160188", X"003f004e",
X"fffe0051", X"00310008", X"ffdbfcd8", X"fe050043", X"ffec0056", X"fefcffb5", X"ffb1001a", X"002fffd9",
X"0326ffbf", X"ffc70021", X"001fffef", X"fff10060", X"00380036", X"03e50260", X"001f002a", X"0045001f",
X"fdfcffac", X"000bffaf", X"0003ffdf", X"fd7e0322", X"ffb60028", X"ffa5ffcf", X"0059fc8a", X"ffee000b",
X"ffe6ffae", X"ffd8ff04", X"ffb1ff9e", X"fcb3ffc4", X"0001ffff", X"0018ffe7", X"ffc90327", X"ffbe000b",
X"0048ffb7", X"02010005", X"01e5ffbc", X"ffaf0046", X"ffaaffed", X"002effb8", X"ffc5ffa8", X"0175ffd7",
X"ffcfffb7", X"01aefd11", X"004a0046", X"fffb02d6", X"0043ffa1", X"02bbfd66", X"0046ffbd", X"0013ffae",
X"004d0168", X"ffbcfc7d", X"fe880042", X"004effb2", X"ff9f0061", X"ffb7ffc6", X"ffc90056", X"ffa5fff7",
X"0005004e", X"000fffda", X"0001027f", X"00420033", X"003bffac", X"feb20008", X"0048ffc9", X"ffa3ffae",
X"014a005c", X"0040ffa2", X"0057fe19", X"fdca0041", X"0018fd62", X"002a000a", X"0026005f", X"fffc016e",
X"ffe3001d", X"ffa2005b", X"fd6c0030", X"0056ffd8", X"03880301", X"ffb4fffc", X"ffd3004e", X"fff2ffb7",
X"ffc6ffba", X"fc97ffbb", X"ffdaff16", X"002effa6", X"ffa3ff9e", X"ffee0025", X"ffd40058", X"0061fdd7",
X"ffc7fe2b", X"ffd6ffc6", X"01720025", X"012bfeb5", X"ffabffcf", X"00b40055", X"012e0396", X"ffb8ff80",
X"ffe6fff5", X"ffe7ffc1", X"00050019", X"fff2ffd1", X"00450038", X"fc1e020d", X"fd870215", X"ffcbffff",
X"fff6ffd2", X"ffcb0062", X"fff3004e", X"ffbe0042", X"ffcf0031", X"ffbefff7", X"03590012", X"ffb80048",
X"000b00bd", X"001dffc7", X"ffcd0051", X"0001fd42", X"ffc2002d", X"fff7ffe3", X"00400036", X"fd13feb6",
X"fff8ffab", X"fecbffaf", X"0052fe7c", X"005cffa8", X"0062ffc6", X"ffcf002b", X"037efc5a", X"ffd1ffa2",
X"fccdffde", X"fca5fd1b", X"005c0006", X"004bffb7", X"fc3b0015", X"0022ffa6", X"fdb400fc", X"fd1effc0",
X"ffbeffa0", X"ffe40042", X"ffbfffed", X"0020ffaa", X"01c90015", X"fe9c0016", X"027b017a", X"ffbd001f",
X"0060004f", X"ffbf025c", X"002f002b", X"ffc4ffbf", X"ffb503cf", X"ffbaffe2", X"ffb7ffcb", X"ffce005b",
X"ffcdfc61", X"0031ffd7", X"0029ffa7", X"fd580003", X"014f033d", X"0015ffac", X"fcfa0229", X"ffa6005a",
X"000bffa6", X"fcf30031", X"005dffae", X"0052010b", X"00160033", X"0061004e", X"03de032d", X"ffde0022",
X"004d0052", X"ffc10045", X"ffabff8e", X"ffb70007", X"fff5001b", X"004f0005", X"000c0058", X"fcd1005f",
X"fc48ffb0", X"fe89fd14", X"003effa9", X"ffebffb1", X"0031ffcf", X"ffd00030", X"fffe0002", X"0006feb8",
X"ff9e0009", X"ffee001d", X"00420023", X"004cffb3", X"ffc6003a", X"000c021c", X"02af0030", X"fc570041",
X"fffefff3", X"ff9efe86", X"fc270039", X"fff7ffe9", X"ffa6ffc0", X"001cfff6", X"ff9f00ac", X"000301c2",
X"00060008", X"005c0058", X"0042003c", X"0052001d", X"002c003b", X"ff9d0030", X"fe8f003c", X"00160058",
X"ffc1ffbe", X"00280059", X"003affe8", X"ff16001a", X"02b00053", X"0057ffdb", X"0037fc25", X"0023ffc9",
X"004e000b", X"ffa1fff4", X"003a0019", X"004d0031", X"fef6004a", X"00630042", X"fcf7000b", X"0036003a",
X"003efff9", X"003b004d", X"0030ffac", X"ffd70029", X"ffbd0044", X"004affe3", X"ffad0036", X"ffa4ffa6",
X"0034ffa9", X"03a6ffe0", X"ffba0039", X"002e0015", X"0034002c", X"ff6dffcc", X"0045005e", X"ffd1ffed",
X"ffa1ffa7", X"0010ffc7", X"005c003c", X"00100048", X"0050002d", X"00f5ffa6", X"007cffbb", X"fff5003a",
X"ffb20047", X"005effd8", X"fff5ffad", X"ffd9ffd5", X"001effce", X"fff9ffca", X"fcff03a4", X"010a0022",
X"feecffb0", X"02f6fffe", X"fd920016", X"0032fd43", X"fff4003f", X"021f003a", X"fffa0063", X"03280006",
X"0066fdb5", X"ffc9ffa1", X"023affde", X"fff0fff7", X"ffec0002", X"001effc1", X"00070043", X"0040ffbb",
X"fffd0062", X"000d0003", X"ff0f0040", X"0044fffc", X"fffaffc2", X"00310044", X"0023ffac", X"0017ffe9",
X"fff1ffab", X"02240034", X"0030ffdd", X"023bffcc", X"ffc5fe50", X"fff5ffd7", X"000a0001", X"ffc4ffb1",
X"ffcf0027", X"000efc4a", X"ffcd005e", X"fd5a002a", X"ffc4ffea", X"004e0052", X"0375ffd7", X"ffc3004a",
X"0027ffe9", X"ffd5ffd4", X"fff7000e", X"ffbbffa5", X"002dffe1", X"004dffb0", X"ffb4ffb8", X"ffb8004e",
X"00710057", X"fd07ffd8", X"005bfff7", X"004e0052", X"01a80029", X"ffd90018", X"fff10009", X"ffac000f",
X"0122fff0", X"ffdb0383", X"004f0036", X"ffc1ffe7", X"ffdcffc3", X"ffbf0037", X"0033ffa2", X"ffec0035",
X"005bffb9", X"ffacfff0", X"0010fce2", X"fff9fff5", X"0215ffa1", X"ffdf0051", X"ffc0ffea", X"fda3fffb",
X"0043000a", X"ffe1ffdc", X"005cfff3", X"005bfe5b", X"01f5ffed", X"0048002b", X"00300006", X"0045001f",
X"0030fff3", X"004c0059", X"ffdfffee", X"ffe8004b", X"ffe00020", X"0335000b", X"0051ffe0", X"01300013",
X"fffe0128", X"ffceff9e", X"ffcdfff5", X"ffe003cc", X"fff10057", X"0286fda7", X"004b0050", X"ffb002a8",
X"0059000b", X"ffab000d", X"0061002a", X"001b0380", X"ffc20047", X"003d00b4", X"02280168", X"00ab0041",
X"ffbc000c", X"001e0044", X"005afcc2", X"ffaf000a", X"ff5dffc8", X"002dffe4", X"0020000b", X"ffd4fff0",
X"fffaff5f", X"0039ffa6", X"ffc5003b", X"fc7fffca", X"0048ffd5", X"00260248", X"0027ffc0", X"03860017",
X"0028004a", X"fccbffa3", X"ffd2002e", X"ffccffc2", X"0038ffaa", X"0047002c", X"005d0150", X"00400097",
X"fdd6ffc3", X"ffdb0032", X"fd90000b", X"ffbc0044", X"0008ffd6", X"fc20ffca", X"027e001c", X"000bfdb7",
X"ffe2fff0", X"ffe5ffbe", X"005c001b", X"002bffa3", X"000c01ca", X"ffab0058", X"fffeffe6", X"008affa9",
X"02aa003e", X"0008ffae", X"000fffd1", X"0007ffc6", X"001b0043", X"00300021", X"fe1bff3e", X"ffd40125",
X"0004001e", X"0035fffc", X"000a0026", X"fff20060", X"fff6ffad", X"0017ffe1", X"0026fff6", X"00580002",
X"00150034", X"010e001b", X"ffa4002a", X"03370049", X"002ffdb2", X"0007ffb1", X"ffe6ffb1", X"fcea0272",
X"ffbdffb7", X"fe46ffce", X"000fffda", X"004affcd", X"ffd20033", X"fff8ff9f", X"0154ffd8", X"003dffc3",
X"ffbfffdd", X"0028fe01", X"003e003a", X"0046ffed", X"ffe5fce2", X"004402ec", X"002d0360", X"0043fe91",
X"003effe7", X"fff3003f", X"fea0ffb5", X"0055ffc2", X"0051ffad", X"ffd70027", X"fffeffb1", X"fef70002",
X"ffccffad", X"fff0ffac", X"01b3ffdc", X"ffba001b", X"0025ffce", X"0047fff2", X"ffa2fffa", X"feb3012e",
X"ffd2001f", X"ffde002e", X"ffa70086", X"005e005f", X"fffe0002", X"005c0008", X"0023016d", X"ffb5ff1f",
X"ffd1fff4", X"0041022f", X"fff00033", X"0018004c", X"0061ffd1", X"ffe40032", X"fffefc87", X"ffc2ffed",
X"fe38ffc1", X"ffa7ffaf", X"001f01e6", X"003002d4", X"001fffb6", X"ffe60045", X"001f012d", X"002a028c",
X"0023fefb", X"004f0032", X"fff900ab", X"fe7e0007", X"001a0056", X"ffd0018b", X"ffeeffc9", X"0017022b",
X"ffdb003b", X"ffc0ffe7", X"0003ffcd", X"ffe30345", X"005b00e5", X"0046fe6a", X"fc2e0063", X"ffedffb4",
X"004e0059", X"0016002f", X"002fffef", X"000d0035", X"00570035", X"feff0004", X"ffc1024a", X"ffc4fe31",
X"005f0005", X"00220042", X"002fff3d", X"00020006", X"ffebffd9", X"002c0038", X"ffc3ffad", X"0223fcfe",
X"ffcb0005", X"0371ffbe", X"02670055", X"fff30013", X"ffd1ff4d", X"ffcb0140", X"005effd7", X"004effa1",
X"0024fccd", X"03c9ffdc", X"ffd4fff7", X"ffdcffa7", X"ffe7fff9", X"00450008", X"ffa2ffd7", X"03620301",
X"0027038b", X"ffef0003", X"0032ffaa", X"ffcdffce", X"0017fd32", X"00320032", X"004600e6", X"ffc4ffa2",
X"0044fc6e", X"0038ffdc", X"0025ffec", X"017effdb", X"037ffff5", X"ffcdffbe", X"ffd90057", X"ffa8fff7",
X"ffcc001b", X"02a0ffe8", X"ffa00005", X"ffa7004a", X"fff403e1", X"0027001c", X"000cfe2f", X"0016001f",
X"ffe0ffbf", X"ffa7fc9f", X"ffdbffb3", X"fff70009", X"fe86ffdb", X"fff2ffab", X"ffd3ffaa", X"0028002d",
X"ffd8ffd8", X"ffa801fb", X"ffabffc5", X"ff9d0041", X"ffe203a1", X"0287ffb5", X"012dffb8", X"ffe80028",
X"0036ffaf", X"ffa3000a", X"0017fffe", X"0291005c", X"0010ffb7", X"feabffb1", X"002dfc53", X"fff2fffc",
X"004bffed", X"0045ffd6", X"ffddffbb", X"fdaf0014", X"fda1ffa3", X"00040008", X"001d00a7", X"ffcc0034",
X"ffde023e", X"00070035", X"00620328", X"002dfe0d", X"ffcc0008", X"ffcc0010", X"032cffb7", X"0012fff5",
X"ffb8003f", X"0003fff7", X"005cfffd", X"fcd70011", X"0038002c", X"ffc3fec2", X"ffa3ffbc", X"000cfff7",
X"0053002e", X"01fe0033", X"0007002f", X"003efecd", X"ffd00056", X"ff22ffb9", X"fff8fffa", X"ffdfffae",
X"ffdb0016", X"fffa002f", X"0056000e", X"00930060", X"fff1ffd1", X"ff9e0042", X"003d004d", X"fceb0062",
X"fc2e0052", X"004ffcdc", X"0061ffb1", X"ffd50387", X"001a02cd", X"ffae0020", X"ffd6fd3c", X"0050fe84",
X"002a0039", X"ffc4003d", X"fffcffa0", X"fff20022", X"fffdfff2", X"003dff35", X"fff0ffd3", X"001d012b",
X"0008ffe4", X"fe9efff5", X"ffeaffb6", X"001cffb5", X"ffa6fff6", X"fff40063", X"ff4d000d", X"ffb70030",
X"ffadffd2", X"fff6002b", X"001b0049", X"ffad0034", X"ffadffbb", X"ff9effb0", X"fff9fe11", X"01beffdb",
X"0044fff2", X"0041ffbf", X"006fffe2", X"ffa10043", X"005b005e", X"005cffac", X"fe15ffd4", X"fffbfff5",
X"00090060", X"ffde0160", X"000d000c", X"ffe1ff9e", X"fffd0056", X"00530003", X"0047ffca", X"ffd502e7",
X"ffbb002c", X"ffa60019", X"ffa001b8", X"0046fdf4", X"03a5ffdf", X"0004fccd", X"0039ffee", X"ff02004c",
X"ffdafff8", X"ffcbffcf", X"ffb4ffdf", X"fc9dffea", X"ffbcffdb", X"fe780005", X"ff9fffd9", X"ffccffb8",
X"fff2fcb0", X"ffa5ffad", X"ffe80058", X"011d0018", X"ffcf0032", X"001c000e", X"025d0055", X"ffa3002f",
X"fff1002b", X"002c0038", X"00530021", X"ffa4000c", X"0051fc44", X"ff0cffc3", X"001f001f", X"000a001b",
X"ffc5ffc9", X"002cfff8", X"0342ffb3", X"00320042", X"0007ffce", X"ffd80021", X"ffdbffd5", X"0008003f",
X"0265ff34", X"036f0015", X"03580020", X"002d000c", X"ff9effee", X"ffcb0018", X"ffcfffae", X"ffc70058",
X"00240002", X"0018ffb0", X"0044ffae", X"0005fcfb", X"fcd1ffe6", X"03c8fd82", X"0343ffe8", X"ffa1ffa3",
X"001b0058", X"004cffe9", X"00180254", X"ffc2003d", X"fffe0001", X"fd9bff9e", X"ffbe0002", X"ffc40025",
X"ffb1ffdd", X"ff0effd1", X"0040005d", X"ffbd005e", X"ffe40013", X"ffdd003f", X"fe50ffad", X"0040ffab",
X"fc990024", X"021effe3", X"fc31ffd6", X"0005ffa8", X"fffdffd3", X"ffed0048", X"004effe7", X"ffcaffa1",
X"00390041", X"ffc8001b", X"002affd4", X"001d001d", X"ffa70025", X"0005003f", X"0029ffb8", X"fff4000f",
X"001b002d", X"0061002b", X"0011fff0", X"0043ffbc", X"000c0015", X"0032fffe", X"0004005c", X"00210038",
X"00020044", X"ffd7ffdc", X"ffedff9d", X"fff70022", X"0014ffaa", X"00200051", X"ffd70015", X"ffeeffed",
X"fff40003", X"002afff3", X"0011001f", X"fffeffe0", X"0029ffd9", X"ffd4ffe7", X"ffe3ffe3", X"002d002b",
X"ffe60022", X"ffe00032", X"0016ffda", X"ffd30013", X"00090029", X"ffe50021", X"fff70010", X"fff8fff6",
X"ffd8fff9", X"ffe9000f", X"ffd6ffd2", X"ffee0021", X"fffeffd3", X"000efff8", X"ffe6fff1", X"ffd9000f",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000"
	);

begin

	-- port A
	process(clka)
	begin
		if rising_edge(clka) then
			if ena = '1' then
				for i in 0 to 3 loop
					if wea(i) = '1' then
						RAM(conv_integer(addra))((i + 1) * 8 - 1 downto i * 8) := dia((i + 1) * 8 - 1 downto i * 8);
					end if;
				end loop;
				doa <= RAM(conv_integer(addra));
			end if;
		end if;
	end process;

	-- port B
	process(clkb)
	begin
		if rising_edge(clkb) then
			if enb = '1' then
				dob <= RAM(conv_integer(addrb));
			end if;
		end if;
	end process;
end rtl;
