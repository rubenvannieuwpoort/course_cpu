library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_types.all;
use work.core_constants.all;


entity decode is
	port (
		clk: in std_logic;
		input: in fetch_output_t;
		output: out decode_output_t := DEFAULT_DECODE_OUTPUT
	);
end decode;


architecture rtl of decode is
begin

	process (clk)
	begin
		if rising_edge(clk) then
			if input.is_active = '1' then
				-- TODO: decode instructions
			else
				output <= DEFAULT_DECODE_OUTPUT;
			end if;
		end if;
	end process;

end rtl;
