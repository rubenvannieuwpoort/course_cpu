library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity decode is
	port (
		clk_in: in std_logic
	);
end decode;


architecture behavioral of decode is
begin
end behavioral;
