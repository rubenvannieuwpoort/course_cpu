library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity top_level is
	port (
		clk_in: in std_logic
	);
end top_level;


architecture rtl of top_level is
begin
end rtl;
