library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity fetch is
	port (
		clk_in: in std_logic
	);
end fetch;


architecture rtl of fetch is
begin
end rtl;
