library ieee;
use ieee.std_logic_1164.all;


package core_types is
	type fetch_output_t is record
	end record fetch_output_t;
end package core_types;
